module aximm();

endmodule
